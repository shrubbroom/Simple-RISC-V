module EX()
